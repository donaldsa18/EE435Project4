/*
* Newspaper FSM states
*
* Authors: Matthew Erhardt, Anthony Donaldson
* Date: 3/23/2018
*
*/
package states;
typedef enum {S0,S5,S10,S15,S20,S25,S30,SHold} state_t;
endpackage
