package prob2states;
typedef enum {S0,S1,S2,S3,S4,S5,S6,S7} state_t;
endpackage