package states;
typedef enum {S0,S5,S10,S15,S20,S25,S30} state_t;
endpackage
